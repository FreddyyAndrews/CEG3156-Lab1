LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY eight_bit_array_multiplier IS 
	PORT
	(
		A :  IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		B :  IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		P :  OUT  STD_LOGIC_VECTOR(17 DOWNTO 0);
		O_first_11 : OUT STD_LOGIC_VECTOR(10 downto 0)
	);
END eight_bit_array_multiplier;

ARCHITECTURE bdf_type OF eight_bit_array_multiplier IS 

COMPONENT array_multiplier_unit
	PORT(a : IN STD_LOGIC	;
		 b : IN STD_LOGIC;
		 c_in : IN STD_LOGIC;
		 pp_in : IN STD_LOGIC;
		 a_through : OUT STD_LOGIC;
		 b_through : OUT STD_LOGIC;
		 c_out : OUT STD_LOGIC;
		 pp_out : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	GND :  STD_LOGIC;
SIGNAL	P_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(17 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_106 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_107 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_108 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_109 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_110 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_111 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_112 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_113 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_114 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_115 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_116 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_117 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_118 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_119 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_120 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_121 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_122 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_123 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_124 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_125 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_126 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_127 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_128 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_129 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_130 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_131 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_132 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_133 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_134 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_135 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_136 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_137 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_138 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_139 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_140 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_141 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_142 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_143 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_144 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_145 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_146 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_147 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_148 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_149 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_150 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_151 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_152 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_153 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_154 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_155 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_156 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_157 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_158 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_159 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_160 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_161 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_162 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_163 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_164 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_165 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_166 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_167 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_168 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_169 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_170 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_171 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_172 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_173 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_174 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_175 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_176 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_177 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_178 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_179 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_180 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_181 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_182 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_183 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_184 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_185 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_186 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_187 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_188 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_189 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_190 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_191 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_192 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_193 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_194 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_195 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_196 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_197 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_198 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_199 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_200 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_201 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_202 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_203 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_204 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_205 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_206 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_207 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_208 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_209 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_210 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_211 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_212 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_213 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_214 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_215 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_216 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_217 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_218 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_219 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_220 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_221 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_222 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_223 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_224 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_225 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_226 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_227 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_228 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_229 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_230 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_231 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_232 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_233 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_234 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_235 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_236 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_237 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_238 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_239 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_240 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_241 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_242 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_243 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_244 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_245 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_246 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_247 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_248 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_249 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_250 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_251 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_252 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_253 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_254 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_255 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_256 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_257 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_258 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_259 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_260 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_261 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_262 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_263 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_264 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_265 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_266 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_267 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_268 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_269 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_270 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_271 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_272 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_273 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_274 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_275 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_276 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_277 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_278 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_279 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_280 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_281 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_282 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_283 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_284 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_285 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_286 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_287 :  STD_LOGIC;


BEGIN 



b2v_inst : array_multiplier_unit
PORT MAP(a => A(0),
		 b => B(0),
		 c_in => GND,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_92,
		 b_through => SYNTHESIZED_WIRE_58,
		 c_out => SYNTHESIZED_WIRE_59,
		 pp_out => P_ALTERA_SYNTHESIZED(0));



b2v_inst100 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_0,
		 b => SYNTHESIZED_WIRE_1,
		 c_in => SYNTHESIZED_WIRE_2,
		 pp_in => SYNTHESIZED_WIRE_3,
		 a_through => SYNTHESIZED_WIRE_4,
		 c_out => SYNTHESIZED_WIRE_7,
		 pp_out => SYNTHESIZED_WIRE_161);


b2v_inst101 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_4,
		 b => SYNTHESIZED_WIRE_5,
		 c_in => SYNTHESIZED_WIRE_6,
		 pp_in => SYNTHESIZED_WIRE_7,
		 a_through => SYNTHESIZED_WIRE_8,
		 c_out => SYNTHESIZED_WIRE_11,
		 pp_out => SYNTHESIZED_WIRE_191);


b2v_inst102 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_8,
		 b => SYNTHESIZED_WIRE_9,
		 c_in => SYNTHESIZED_WIRE_10,
		 pp_in => SYNTHESIZED_WIRE_11,
		 a_through => SYNTHESIZED_WIRE_12,
		 c_out => SYNTHESIZED_WIRE_15,
		 pp_out => SYNTHESIZED_WIRE_221);


b2v_inst103 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_12,
		 b => SYNTHESIZED_WIRE_13,
		 c_in => SYNTHESIZED_WIRE_14,
		 pp_in => SYNTHESIZED_WIRE_15,
		 a_through => SYNTHESIZED_WIRE_16,
		 c_out => SYNTHESIZED_WIRE_19,
		 pp_out => SYNTHESIZED_WIRE_251);


b2v_inst104 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_16,
		 b => SYNTHESIZED_WIRE_17,
		 c_in => SYNTHESIZED_WIRE_18,
		 pp_in => SYNTHESIZED_WIRE_19,
		 a_through => SYNTHESIZED_WIRE_50,
		 c_out => SYNTHESIZED_WIRE_53,
		 pp_out => SYNTHESIZED_WIRE_281);


b2v_inst105 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_20,
		 b => B(8),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_21,
		 b_through => SYNTHESIZED_WIRE_23,
		 c_out => SYNTHESIZED_WIRE_24,
		 pp_out => P_ALTERA_SYNTHESIZED(8));


b2v_inst106 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_22,
		 b => SYNTHESIZED_WIRE_23,
		 c_in => SYNTHESIZED_WIRE_24,
		 pp_in => SYNTHESIZED_WIRE_25,
		 b_through => SYNTHESIZED_WIRE_27,
		 c_out => SYNTHESIZED_WIRE_28,
		 pp_out => P_ALTERA_SYNTHESIZED(9));


b2v_inst107 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_26,
		 b => SYNTHESIZED_WIRE_27,
		 c_in => SYNTHESIZED_WIRE_28,
		 pp_in => SYNTHESIZED_WIRE_29,
		 b_through => SYNTHESIZED_WIRE_31,
		 c_out => SYNTHESIZED_WIRE_32,
		 pp_out => P_ALTERA_SYNTHESIZED(10));


b2v_inst108 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_30,
		 b => SYNTHESIZED_WIRE_31,
		 c_in => SYNTHESIZED_WIRE_32,
		 pp_in => SYNTHESIZED_WIRE_33,
		 b_through => SYNTHESIZED_WIRE_35,
		 c_out => SYNTHESIZED_WIRE_36,
		 pp_out => P_ALTERA_SYNTHESIZED(11));


b2v_inst109 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_34,
		 b => SYNTHESIZED_WIRE_35,
		 c_in => SYNTHESIZED_WIRE_36,
		 pp_in => SYNTHESIZED_WIRE_37,
		 b_through => SYNTHESIZED_WIRE_39,
		 c_out => SYNTHESIZED_WIRE_40,
		 pp_out => P_ALTERA_SYNTHESIZED(12));


b2v_inst110 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_38,
		 b => SYNTHESIZED_WIRE_39,
		 c_in => SYNTHESIZED_WIRE_40,
		 pp_in => SYNTHESIZED_WIRE_41,
		 b_through => SYNTHESIZED_WIRE_43,
		 c_out => SYNTHESIZED_WIRE_44,
		 pp_out => P_ALTERA_SYNTHESIZED(13));


b2v_inst111 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_42,
		 b => SYNTHESIZED_WIRE_43,
		 c_in => SYNTHESIZED_WIRE_44,
		 pp_in => SYNTHESIZED_WIRE_45,
		 b_through => SYNTHESIZED_WIRE_47,
		 c_out => SYNTHESIZED_WIRE_48,
		 pp_out => P_ALTERA_SYNTHESIZED(14));


b2v_inst112 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_46,
		 b => SYNTHESIZED_WIRE_47,
		 c_in => SYNTHESIZED_WIRE_48,
		 pp_in => SYNTHESIZED_WIRE_49,
		 b_through => SYNTHESIZED_WIRE_55,
		 c_out => SYNTHESIZED_WIRE_56,
		 pp_out => P_ALTERA_SYNTHESIZED(15));


b2v_inst113 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_50,
		 b => SYNTHESIZED_WIRE_51,
		 c_in => SYNTHESIZED_WIRE_52,
		 pp_in => SYNTHESIZED_WIRE_53,
		 a_through => SYNTHESIZED_WIRE_54,
		 c_out => SYNTHESIZED_WIRE_57,
		 pp_out => SYNTHESIZED_WIRE_49);


b2v_inst114 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_54,
		 b => SYNTHESIZED_WIRE_55,
		 c_in => SYNTHESIZED_WIRE_56,
		 pp_in => SYNTHESIZED_WIRE_57,
		 c_out => P_ALTERA_SYNTHESIZED(17),
		 pp_out => P_ALTERA_SYNTHESIZED(16));


b2v_inst35 : array_multiplier_unit
PORT MAP(a => A(1),
		 b => SYNTHESIZED_WIRE_58,
		 c_in => SYNTHESIZED_WIRE_59,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_66,
		 b_through => SYNTHESIZED_WIRE_86,
		 c_out => SYNTHESIZED_WIRE_87,
		 pp_out => SYNTHESIZED_WIRE_93);


b2v_inst36 : array_multiplier_unit
PORT MAP(a => A(3),
		 b => SYNTHESIZED_WIRE_60,
		 c_in => SYNTHESIZED_WIRE_61,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_70,
		 b_through => SYNTHESIZED_WIRE_88,
		 c_out => SYNTHESIZED_WIRE_89,
		 pp_out => SYNTHESIZED_WIRE_97);


b2v_inst37 : array_multiplier_unit
PORT MAP(a => A(5),
		 b => SYNTHESIZED_WIRE_62,
		 c_in => SYNTHESIZED_WIRE_63,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_74,
		 b_through => SYNTHESIZED_WIRE_90,
		 c_out => SYNTHESIZED_WIRE_91,
		 pp_out => SYNTHESIZED_WIRE_101);


b2v_inst38 : array_multiplier_unit
PORT MAP(a => A(7),
		 b => SYNTHESIZED_WIRE_64,
		 c_in => SYNTHESIZED_WIRE_65,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_78,
		 b_through => SYNTHESIZED_WIRE_282,
		 c_out => SYNTHESIZED_WIRE_283,
		 pp_out => SYNTHESIZED_WIRE_105);


b2v_inst39 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_66,
		 b => SYNTHESIZED_WIRE_67,
		 c_in => SYNTHESIZED_WIRE_68,
		 pp_in => SYNTHESIZED_WIRE_69,
		 a_through => SYNTHESIZED_WIRE_82,
		 b_through => SYNTHESIZED_WIRE_95,
		 c_out => SYNTHESIZED_WIRE_96,
		 pp_out => SYNTHESIZED_WIRE_107);


b2v_inst40 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_70,
		 b => SYNTHESIZED_WIRE_71,
		 c_in => SYNTHESIZED_WIRE_72,
		 pp_in => SYNTHESIZED_WIRE_73,
		 a_through => SYNTHESIZED_WIRE_112,
		 b_through => SYNTHESIZED_WIRE_99,
		 c_out => SYNTHESIZED_WIRE_100,
		 pp_out => SYNTHESIZED_WIRE_111);


b2v_inst41 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_74,
		 b => SYNTHESIZED_WIRE_75,
		 c_in => SYNTHESIZED_WIRE_76,
		 pp_in => SYNTHESIZED_WIRE_77,
		 a_through => SYNTHESIZED_WIRE_120,
		 b_through => SYNTHESIZED_WIRE_103,
		 c_out => SYNTHESIZED_WIRE_104,
		 pp_out => SYNTHESIZED_WIRE_119);


b2v_inst42 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_78,
		 b => SYNTHESIZED_WIRE_79,
		 c_in => SYNTHESIZED_WIRE_80,
		 pp_in => SYNTHESIZED_WIRE_81,
		 a_through => SYNTHESIZED_WIRE_128,
		 b_through => SYNTHESIZED_WIRE_285,
		 c_out => SYNTHESIZED_WIRE_286,
		 pp_out => SYNTHESIZED_WIRE_127);


b2v_inst43 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_82,
		 b => SYNTHESIZED_WIRE_83,
		 c_in => SYNTHESIZED_WIRE_84,
		 pp_in => SYNTHESIZED_WIRE_85,
		 a_through => SYNTHESIZED_WIRE_134,
		 b_through => SYNTHESIZED_WIRE_109,
		 c_out => SYNTHESIZED_WIRE_110,
		 pp_out => SYNTHESIZED_WIRE_133);


b2v_inst44 : array_multiplier_unit
PORT MAP(a => A(2),
		 b => SYNTHESIZED_WIRE_86,
		 c_in => SYNTHESIZED_WIRE_87,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_94,
		 b_through => SYNTHESIZED_WIRE_60,
		 c_out => SYNTHESIZED_WIRE_61,
		 pp_out => SYNTHESIZED_WIRE_69);


b2v_inst45 : array_multiplier_unit
PORT MAP(a => A(4),
		 b => SYNTHESIZED_WIRE_88,
		 c_in => SYNTHESIZED_WIRE_89,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_98,
		 b_through => SYNTHESIZED_WIRE_62,
		 c_out => SYNTHESIZED_WIRE_63,
		 pp_out => SYNTHESIZED_WIRE_73);


b2v_inst46 : array_multiplier_unit
PORT MAP(a => A(6),
		 b => SYNTHESIZED_WIRE_90,
		 c_in => SYNTHESIZED_WIRE_91,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_102,
		 b_through => SYNTHESIZED_WIRE_64,
		 c_out => SYNTHESIZED_WIRE_65,
		 pp_out => SYNTHESIZED_WIRE_77);


b2v_inst47 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_92,
		 b => B(1),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_93,
		 a_through => SYNTHESIZED_WIRE_106,
		 b_through => SYNTHESIZED_WIRE_67,
		 c_out => SYNTHESIZED_WIRE_68,
		 pp_out => P_ALTERA_SYNTHESIZED(1));


b2v_inst48 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_94,
		 b => SYNTHESIZED_WIRE_95,
		 c_in => SYNTHESIZED_WIRE_96,
		 pp_in => SYNTHESIZED_WIRE_97,
		 a_through => SYNTHESIZED_WIRE_108,
		 b_through => SYNTHESIZED_WIRE_71,
		 c_out => SYNTHESIZED_WIRE_72,
		 pp_out => SYNTHESIZED_WIRE_85);


b2v_inst49 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_98,
		 b => SYNTHESIZED_WIRE_99,
		 c_in => SYNTHESIZED_WIRE_100,
		 pp_in => SYNTHESIZED_WIRE_101,
		 a_through => SYNTHESIZED_WIRE_116,
		 b_through => SYNTHESIZED_WIRE_75,
		 c_out => SYNTHESIZED_WIRE_76,
		 pp_out => SYNTHESIZED_WIRE_115);


b2v_inst50 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_102,
		 b => SYNTHESIZED_WIRE_103,
		 c_in => SYNTHESIZED_WIRE_104,
		 pp_in => SYNTHESIZED_WIRE_105,
		 a_through => SYNTHESIZED_WIRE_124,
		 b_through => SYNTHESIZED_WIRE_79,
		 c_out => SYNTHESIZED_WIRE_80,
		 pp_out => SYNTHESIZED_WIRE_123);


b2v_inst51 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_106,
		 b => B(2),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_107,
		 a_through => SYNTHESIZED_WIRE_132,
		 b_through => SYNTHESIZED_WIRE_83,
		 c_out => SYNTHESIZED_WIRE_84,
		 pp_out => P_ALTERA_SYNTHESIZED(2));


b2v_inst52 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_108,
		 b => SYNTHESIZED_WIRE_109,
		 c_in => SYNTHESIZED_WIRE_110,
		 pp_in => SYNTHESIZED_WIRE_111,
		 a_through => SYNTHESIZED_WIRE_138,
		 b_through => SYNTHESIZED_WIRE_113,
		 c_out => SYNTHESIZED_WIRE_114,
		 pp_out => SYNTHESIZED_WIRE_137);


b2v_inst53 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_112,
		 b => SYNTHESIZED_WIRE_113,
		 c_in => SYNTHESIZED_WIRE_114,
		 pp_in => SYNTHESIZED_WIRE_115,
		 a_through => SYNTHESIZED_WIRE_142,
		 b_through => SYNTHESIZED_WIRE_117,
		 c_out => SYNTHESIZED_WIRE_118,
		 pp_out => SYNTHESIZED_WIRE_141);


b2v_inst54 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_116,
		 b => SYNTHESIZED_WIRE_117,
		 c_in => SYNTHESIZED_WIRE_118,
		 pp_in => SYNTHESIZED_WIRE_119,
		 a_through => SYNTHESIZED_WIRE_146,
		 b_through => SYNTHESIZED_WIRE_121,
		 c_out => SYNTHESIZED_WIRE_122,
		 pp_out => SYNTHESIZED_WIRE_145);


b2v_inst55 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_120,
		 b => SYNTHESIZED_WIRE_121,
		 c_in => SYNTHESIZED_WIRE_122,
		 pp_in => SYNTHESIZED_WIRE_123,
		 a_through => SYNTHESIZED_WIRE_150,
		 b_through => SYNTHESIZED_WIRE_125,
		 c_out => SYNTHESIZED_WIRE_126,
		 pp_out => SYNTHESIZED_WIRE_149);


b2v_inst56 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_124,
		 b => SYNTHESIZED_WIRE_125,
		 c_in => SYNTHESIZED_WIRE_126,
		 pp_in => SYNTHESIZED_WIRE_127,
		 a_through => SYNTHESIZED_WIRE_154,
		 b_through => SYNTHESIZED_WIRE_129,
		 c_out => SYNTHESIZED_WIRE_130,
		 pp_out => SYNTHESIZED_WIRE_153);


b2v_inst57 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_128,
		 b => SYNTHESIZED_WIRE_129,
		 c_in => SYNTHESIZED_WIRE_130,
		 pp_in => SYNTHESIZED_WIRE_131,
		 a_through => SYNTHESIZED_WIRE_158,
		 b_through => SYNTHESIZED_WIRE_1,
		 c_out => SYNTHESIZED_WIRE_2,
		 pp_out => SYNTHESIZED_WIRE_157);


b2v_inst58 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_132,
		 b => B(3),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_133,
		 a_through => SYNTHESIZED_WIRE_162,
		 b_through => SYNTHESIZED_WIRE_135,
		 c_out => SYNTHESIZED_WIRE_136,
		 pp_out => P_ALTERA_SYNTHESIZED(3));


b2v_inst59 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_134,
		 b => SYNTHESIZED_WIRE_135,
		 c_in => SYNTHESIZED_WIRE_136,
		 pp_in => SYNTHESIZED_WIRE_137,
		 a_through => SYNTHESIZED_WIRE_164,
		 b_through => SYNTHESIZED_WIRE_139,
		 c_out => SYNTHESIZED_WIRE_140,
		 pp_out => SYNTHESIZED_WIRE_163);


b2v_inst60 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_138,
		 b => SYNTHESIZED_WIRE_139,
		 c_in => SYNTHESIZED_WIRE_140,
		 pp_in => SYNTHESIZED_WIRE_141,
		 a_through => SYNTHESIZED_WIRE_168,
		 b_through => SYNTHESIZED_WIRE_143,
		 c_out => SYNTHESIZED_WIRE_144,
		 pp_out => SYNTHESIZED_WIRE_167);


b2v_inst61 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_142,
		 b => SYNTHESIZED_WIRE_143,
		 c_in => SYNTHESIZED_WIRE_144,
		 pp_in => SYNTHESIZED_WIRE_145,
		 a_through => SYNTHESIZED_WIRE_172,
		 b_through => SYNTHESIZED_WIRE_147,
		 c_out => SYNTHESIZED_WIRE_148,
		 pp_out => SYNTHESIZED_WIRE_171);


b2v_inst62 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_146,
		 b => SYNTHESIZED_WIRE_147,
		 c_in => SYNTHESIZED_WIRE_148,
		 pp_in => SYNTHESIZED_WIRE_149,
		 a_through => SYNTHESIZED_WIRE_176,
		 b_through => SYNTHESIZED_WIRE_151,
		 c_out => SYNTHESIZED_WIRE_152,
		 pp_out => SYNTHESIZED_WIRE_175);


b2v_inst63 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_150,
		 b => SYNTHESIZED_WIRE_151,
		 c_in => SYNTHESIZED_WIRE_152,
		 pp_in => SYNTHESIZED_WIRE_153,
		 a_through => SYNTHESIZED_WIRE_180,
		 b_through => SYNTHESIZED_WIRE_155,
		 c_out => SYNTHESIZED_WIRE_156,
		 pp_out => SYNTHESIZED_WIRE_179);


b2v_inst64 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_154,
		 b => SYNTHESIZED_WIRE_155,
		 c_in => SYNTHESIZED_WIRE_156,
		 pp_in => SYNTHESIZED_WIRE_157,
		 a_through => SYNTHESIZED_WIRE_184,
		 b_through => SYNTHESIZED_WIRE_159,
		 c_out => SYNTHESIZED_WIRE_160,
		 pp_out => SYNTHESIZED_WIRE_183);


b2v_inst65 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_158,
		 b => SYNTHESIZED_WIRE_159,
		 c_in => SYNTHESIZED_WIRE_160,
		 pp_in => SYNTHESIZED_WIRE_161,
		 a_through => SYNTHESIZED_WIRE_188,
		 b_through => SYNTHESIZED_WIRE_5,
		 c_out => SYNTHESIZED_WIRE_6,
		 pp_out => SYNTHESIZED_WIRE_187);


b2v_inst66 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_162,
		 b => B(4),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_163,
		 a_through => SYNTHESIZED_WIRE_192,
		 b_through => SYNTHESIZED_WIRE_165,
		 c_out => SYNTHESIZED_WIRE_166,
		 pp_out => P_ALTERA_SYNTHESIZED(4));


b2v_inst67 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_164,
		 b => SYNTHESIZED_WIRE_165,
		 c_in => SYNTHESIZED_WIRE_166,
		 pp_in => SYNTHESIZED_WIRE_167,
		 a_through => SYNTHESIZED_WIRE_194,
		 b_through => SYNTHESIZED_WIRE_169,
		 c_out => SYNTHESIZED_WIRE_170,
		 pp_out => SYNTHESIZED_WIRE_193);


b2v_inst68 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_168,
		 b => SYNTHESIZED_WIRE_169,
		 c_in => SYNTHESIZED_WIRE_170,
		 pp_in => SYNTHESIZED_WIRE_171,
		 a_through => SYNTHESIZED_WIRE_198,
		 b_through => SYNTHESIZED_WIRE_173,
		 c_out => SYNTHESIZED_WIRE_174,
		 pp_out => SYNTHESIZED_WIRE_197);


b2v_inst69 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_172,
		 b => SYNTHESIZED_WIRE_173,
		 c_in => SYNTHESIZED_WIRE_174,
		 pp_in => SYNTHESIZED_WIRE_175,
		 a_through => SYNTHESIZED_WIRE_202,
		 b_through => SYNTHESIZED_WIRE_177,
		 c_out => SYNTHESIZED_WIRE_178,
		 pp_out => SYNTHESIZED_WIRE_201);


b2v_inst70 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_176,
		 b => SYNTHESIZED_WIRE_177,
		 c_in => SYNTHESIZED_WIRE_178,
		 pp_in => SYNTHESIZED_WIRE_179,
		 a_through => SYNTHESIZED_WIRE_206,
		 b_through => SYNTHESIZED_WIRE_181,
		 c_out => SYNTHESIZED_WIRE_182,
		 pp_out => SYNTHESIZED_WIRE_205);


b2v_inst71 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_180,
		 b => SYNTHESIZED_WIRE_181,
		 c_in => SYNTHESIZED_WIRE_182,
		 pp_in => SYNTHESIZED_WIRE_183,
		 a_through => SYNTHESIZED_WIRE_210,
		 b_through => SYNTHESIZED_WIRE_185,
		 c_out => SYNTHESIZED_WIRE_186,
		 pp_out => SYNTHESIZED_WIRE_209);


b2v_inst72 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_184,
		 b => SYNTHESIZED_WIRE_185,
		 c_in => SYNTHESIZED_WIRE_186,
		 pp_in => SYNTHESIZED_WIRE_187,
		 a_through => SYNTHESIZED_WIRE_214,
		 b_through => SYNTHESIZED_WIRE_189,
		 c_out => SYNTHESIZED_WIRE_190,
		 pp_out => SYNTHESIZED_WIRE_213);


b2v_inst73 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_188,
		 b => SYNTHESIZED_WIRE_189,
		 c_in => SYNTHESIZED_WIRE_190,
		 pp_in => SYNTHESIZED_WIRE_191,
		 a_through => SYNTHESIZED_WIRE_218,
		 b_through => SYNTHESIZED_WIRE_9,
		 c_out => SYNTHESIZED_WIRE_10,
		 pp_out => SYNTHESIZED_WIRE_217);


b2v_inst74 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_192,
		 b => B(5),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_193,
		 a_through => SYNTHESIZED_WIRE_222,
		 b_through => SYNTHESIZED_WIRE_195,
		 c_out => SYNTHESIZED_WIRE_196,
		 pp_out => P_ALTERA_SYNTHESIZED(5));


b2v_inst75 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_194,
		 b => SYNTHESIZED_WIRE_195,
		 c_in => SYNTHESIZED_WIRE_196,
		 pp_in => SYNTHESIZED_WIRE_197,
		 a_through => SYNTHESIZED_WIRE_224,
		 b_through => SYNTHESIZED_WIRE_199,
		 c_out => SYNTHESIZED_WIRE_200,
		 pp_out => SYNTHESIZED_WIRE_223);


b2v_inst76 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_198,
		 b => SYNTHESIZED_WIRE_199,
		 c_in => SYNTHESIZED_WIRE_200,
		 pp_in => SYNTHESIZED_WIRE_201,
		 a_through => SYNTHESIZED_WIRE_228,
		 b_through => SYNTHESIZED_WIRE_203,
		 c_out => SYNTHESIZED_WIRE_204,
		 pp_out => SYNTHESIZED_WIRE_227);


b2v_inst77 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_202,
		 b => SYNTHESIZED_WIRE_203,
		 c_in => SYNTHESIZED_WIRE_204,
		 pp_in => SYNTHESIZED_WIRE_205,
		 a_through => SYNTHESIZED_WIRE_232,
		 b_through => SYNTHESIZED_WIRE_207,
		 c_out => SYNTHESIZED_WIRE_208,
		 pp_out => SYNTHESIZED_WIRE_231);


b2v_inst78 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_206,
		 b => SYNTHESIZED_WIRE_207,
		 c_in => SYNTHESIZED_WIRE_208,
		 pp_in => SYNTHESIZED_WIRE_209,
		 a_through => SYNTHESIZED_WIRE_236,
		 b_through => SYNTHESIZED_WIRE_211,
		 c_out => SYNTHESIZED_WIRE_212,
		 pp_out => SYNTHESIZED_WIRE_235);


b2v_inst79 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_210,
		 b => SYNTHESIZED_WIRE_211,
		 c_in => SYNTHESIZED_WIRE_212,
		 pp_in => SYNTHESIZED_WIRE_213,
		 a_through => SYNTHESIZED_WIRE_240,
		 b_through => SYNTHESIZED_WIRE_215,
		 c_out => SYNTHESIZED_WIRE_216,
		 pp_out => SYNTHESIZED_WIRE_239);


b2v_inst80 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_214,
		 b => SYNTHESIZED_WIRE_215,
		 c_in => SYNTHESIZED_WIRE_216,
		 pp_in => SYNTHESIZED_WIRE_217,
		 a_through => SYNTHESIZED_WIRE_244,
		 b_through => SYNTHESIZED_WIRE_219,
		 c_out => SYNTHESIZED_WIRE_220,
		 pp_out => SYNTHESIZED_WIRE_243);


b2v_inst81 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_218,
		 b => SYNTHESIZED_WIRE_219,
		 c_in => SYNTHESIZED_WIRE_220,
		 pp_in => SYNTHESIZED_WIRE_221,
		 a_through => SYNTHESIZED_WIRE_248,
		 b_through => SYNTHESIZED_WIRE_13,
		 c_out => SYNTHESIZED_WIRE_14,
		 pp_out => SYNTHESIZED_WIRE_247);


b2v_inst82 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_222,
		 b => B(6),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_223,
		 a_through => SYNTHESIZED_WIRE_252,
		 b_through => SYNTHESIZED_WIRE_225,
		 c_out => SYNTHESIZED_WIRE_226,
		 pp_out => P_ALTERA_SYNTHESIZED(6));


b2v_inst83 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_224,
		 b => SYNTHESIZED_WIRE_225,
		 c_in => SYNTHESIZED_WIRE_226,
		 pp_in => SYNTHESIZED_WIRE_227,
		 a_through => SYNTHESIZED_WIRE_254,
		 b_through => SYNTHESIZED_WIRE_229,
		 c_out => SYNTHESIZED_WIRE_230,
		 pp_out => SYNTHESIZED_WIRE_253);


b2v_inst84 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_228,
		 b => SYNTHESIZED_WIRE_229,
		 c_in => SYNTHESIZED_WIRE_230,
		 pp_in => SYNTHESIZED_WIRE_231,
		 a_through => SYNTHESIZED_WIRE_258,
		 b_through => SYNTHESIZED_WIRE_233,
		 c_out => SYNTHESIZED_WIRE_234,
		 pp_out => SYNTHESIZED_WIRE_257);


b2v_inst85 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_232,
		 b => SYNTHESIZED_WIRE_233,
		 c_in => SYNTHESIZED_WIRE_234,
		 pp_in => SYNTHESIZED_WIRE_235,
		 a_through => SYNTHESIZED_WIRE_262,
		 b_through => SYNTHESIZED_WIRE_237,
		 c_out => SYNTHESIZED_WIRE_238,
		 pp_out => SYNTHESIZED_WIRE_261);


b2v_inst86 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_236,
		 b => SYNTHESIZED_WIRE_237,
		 c_in => SYNTHESIZED_WIRE_238,
		 pp_in => SYNTHESIZED_WIRE_239,
		 a_through => SYNTHESIZED_WIRE_266,
		 b_through => SYNTHESIZED_WIRE_241,
		 c_out => SYNTHESIZED_WIRE_242,
		 pp_out => SYNTHESIZED_WIRE_265);


b2v_inst87 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_240,
		 b => SYNTHESIZED_WIRE_241,
		 c_in => SYNTHESIZED_WIRE_242,
		 pp_in => SYNTHESIZED_WIRE_243,
		 a_through => SYNTHESIZED_WIRE_270,
		 b_through => SYNTHESIZED_WIRE_245,
		 c_out => SYNTHESIZED_WIRE_246,
		 pp_out => SYNTHESIZED_WIRE_269);


b2v_inst88 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_244,
		 b => SYNTHESIZED_WIRE_245,
		 c_in => SYNTHESIZED_WIRE_246,
		 pp_in => SYNTHESIZED_WIRE_247,
		 a_through => SYNTHESIZED_WIRE_274,
		 b_through => SYNTHESIZED_WIRE_249,
		 c_out => SYNTHESIZED_WIRE_250,
		 pp_out => SYNTHESIZED_WIRE_273);


b2v_inst89 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_248,
		 b => SYNTHESIZED_WIRE_249,
		 c_in => SYNTHESIZED_WIRE_250,
		 pp_in => SYNTHESIZED_WIRE_251,
		 a_through => SYNTHESIZED_WIRE_278,
		 b_through => SYNTHESIZED_WIRE_17,
		 c_out => SYNTHESIZED_WIRE_18,
		 pp_out => SYNTHESIZED_WIRE_277);


b2v_inst90 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_252,
		 b => B(7),
		 c_in => GND,
		 pp_in => SYNTHESIZED_WIRE_253,
		 a_through => SYNTHESIZED_WIRE_20,
		 b_through => SYNTHESIZED_WIRE_255,
		 c_out => SYNTHESIZED_WIRE_256,
		 pp_out => P_ALTERA_SYNTHESIZED(7));


b2v_inst91 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_254,
		 b => SYNTHESIZED_WIRE_255,
		 c_in => SYNTHESIZED_WIRE_256,
		 pp_in => SYNTHESIZED_WIRE_257,
		 a_through => SYNTHESIZED_WIRE_22,
		 b_through => SYNTHESIZED_WIRE_259,
		 c_out => SYNTHESIZED_WIRE_260,
		 pp_out => SYNTHESIZED_WIRE_21);


b2v_inst92 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_258,
		 b => SYNTHESIZED_WIRE_259,
		 c_in => SYNTHESIZED_WIRE_260,
		 pp_in => SYNTHESIZED_WIRE_261,
		 a_through => SYNTHESIZED_WIRE_26,
		 b_through => SYNTHESIZED_WIRE_263,
		 c_out => SYNTHESIZED_WIRE_264,
		 pp_out => SYNTHESIZED_WIRE_25);


b2v_inst93 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_262,
		 b => SYNTHESIZED_WIRE_263,
		 c_in => SYNTHESIZED_WIRE_264,
		 pp_in => SYNTHESIZED_WIRE_265,
		 a_through => SYNTHESIZED_WIRE_30,
		 b_through => SYNTHESIZED_WIRE_267,
		 c_out => SYNTHESIZED_WIRE_268,
		 pp_out => SYNTHESIZED_WIRE_29);


b2v_inst94 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_266,
		 b => SYNTHESIZED_WIRE_267,
		 c_in => SYNTHESIZED_WIRE_268,
		 pp_in => SYNTHESIZED_WIRE_269,
		 a_through => SYNTHESIZED_WIRE_34,
		 b_through => SYNTHESIZED_WIRE_271,
		 c_out => SYNTHESIZED_WIRE_272,
		 pp_out => SYNTHESIZED_WIRE_33);


b2v_inst95 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_270,
		 b => SYNTHESIZED_WIRE_271,
		 c_in => SYNTHESIZED_WIRE_272,
		 pp_in => SYNTHESIZED_WIRE_273,
		 a_through => SYNTHESIZED_WIRE_38,
		 b_through => SYNTHESIZED_WIRE_275,
		 c_out => SYNTHESIZED_WIRE_276,
		 pp_out => SYNTHESIZED_WIRE_37);


b2v_inst96 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_274,
		 b => SYNTHESIZED_WIRE_275,
		 c_in => SYNTHESIZED_WIRE_276,
		 pp_in => SYNTHESIZED_WIRE_277,
		 a_through => SYNTHESIZED_WIRE_42,
		 b_through => SYNTHESIZED_WIRE_279,
		 c_out => SYNTHESIZED_WIRE_280,
		 pp_out => SYNTHESIZED_WIRE_41);


b2v_inst97 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_278,
		 b => SYNTHESIZED_WIRE_279,
		 c_in => SYNTHESIZED_WIRE_280,
		 pp_in => SYNTHESIZED_WIRE_281,
		 a_through => SYNTHESIZED_WIRE_46,
		 b_through => SYNTHESIZED_WIRE_51,
		 c_out => SYNTHESIZED_WIRE_52,
		 pp_out => SYNTHESIZED_WIRE_45);


b2v_inst98 : array_multiplier_unit
PORT MAP(a => A(8),
		 b => SYNTHESIZED_WIRE_282,
		 c_in => SYNTHESIZED_WIRE_283,
		 pp_in => GND,
		 a_through => SYNTHESIZED_WIRE_284,
		 c_out => SYNTHESIZED_WIRE_287,
		 pp_out => SYNTHESIZED_WIRE_81);


b2v_inst99 : array_multiplier_unit
PORT MAP(a => SYNTHESIZED_WIRE_284,
		 b => SYNTHESIZED_WIRE_285,
		 c_in => SYNTHESIZED_WIRE_286,
		 pp_in => SYNTHESIZED_WIRE_287,
		 a_through => SYNTHESIZED_WIRE_0,
		 c_out => SYNTHESIZED_WIRE_3,
		 pp_out => SYNTHESIZED_WIRE_131);

P <= P_ALTERA_SYNTHESIZED;
O_first_11 <= P_ALTERA_SYNTHESIZED(17 downto 7);

GND <= '0';
END bdf_type;