-- TODO: Implement this file